module Adder (
    in1,
    in2,
    out
);


endmoudle
